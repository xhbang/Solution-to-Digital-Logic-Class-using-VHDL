LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux21 IS
	PORT	(a,b: IN STD_LOGIC;
			   s: IN STD_LOGIC;
			   y: OUT STD_LOGIC);
END ENTITY mux21;

ARCHITECTURE one OF mux21 IS
	BEGIN
		y<=a WHEN s='0' ELSE
		b WHEN s='1';
END ARCHITECTURE one;